
module Xor_M

(
	//Input
	input A,
	input B,
	
	//Output
	output C

);

assign C = A^B;

endmodule
